library ieee;
use ieee.std_logic_1164.all;

-- Prototype and constant declarations
package CommonTypes is
	
	constant BUTTON_ACTIVE: std_logic := '0';
	

end package;



-- Any function declarations
package body CommonTypes is

end package body;

