library ieee;
use ieee.std_logic_1164.all;


package CommonTypes is 
	constant RESET_ACTIVE: std_logic := '0';
end package;



package body CommonTypes is

end package body;
