library ieee;
use ieee.std_logic_1164.ALL;



package LED is 





end package;
